BZh91AY&SY*�LO �_�Px��g߰����P�wd3rh+@%Q�MOL��F��I����2��i��1OSP���   	L�i�F��     � �0�M0  �4�0� �24�<�b~��ꆁ��1���/���"IQ ,@�I�~�6ؗ��י��B�ib��
�k��a���]��B���vC�	D��I��k�����Ak8hv&�?q���C�,3J���6���L�_�X2�J�� 0��Lyʜ�i�/-����q4e׶K8�3!�a��x�L�\P9L�P�8ʐK��0�����P�H=֞$��U�"��0�(K�
4�!z\�Ҋ���X%E��`\9m�u���o7��_�b$H$ؒH �{�#y���u&�R1V�+n�����ʑk�F��d�R&�)@k�p�����\p{��l��(���U��Kl���}K	�����-�,#8�a$�u���O�c|S���s����W�q�c.H喔��{7 �E@/F"0"L����h�)���<�7��%���ݰ�&�mb���j�ƫ�����h'2)J�^'v*�f�haY���P��P5�(�ꆶ{��.e��}�&���Y�M�½��~��1�����.�(�gݒ`��B�$�s�O�lБ�Ω�A�鞅��#�#�fB��ˌ��l|�%h�=8&X%���Y�P.�No�5�^rJ�УѪs��RĐD �����+Z��M@qz&�s" �CU:�H!Lg��C�fhB�	�b����x�F'��=L% *�^��P���Ǳ[1��1��]�a"�$�#������"��!�c�q�q��2٧��d���F4�RT	�M�4-�m��0�E}�X�<�MrAvx���^���+�Zi�n��:`��6�Y�������U����)�Wbx